module ascii_to_utf8();
endmodule : ascii_to_utf8
